module pipeline1
(
 //input[7:0] OPCODE,
 input[15:0] OPCODE,
 //input[4:0] Ri,
 //input[4:0] Rj,
 output reg [3:0] ALUC,
 output reg [1:0] SH,
 output reg KMux,
 output reg MR,
 output reg MW,
 output reg [4:0] Sel_A,
 output reg [5:0] Sel_B,
 output reg [5:0] Sel_C,
 output reg [6:0] Type,
 output reg [9:0] Dadd
 );
	 
			

endmodule
