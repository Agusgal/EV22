module UC2
(
input [4:0]SelA2,
input [5:0]SelB2,
input [8:0]Type2,
input [8:0]Type3,
input [5:0]SelC3,
input [8:0]Type4,
input [5:0]SelC4,
input [8:0]Type5,
input [5:0]SelC5,
output reg HOLD
 );

 
 //Condiciones para Hold: 




 
always @(*)begin


end

endmodule
